/*
 *		C言語で記述されたアプリケーションから，TECSベースのタイマドラ
 *		イバシミュレータ制御を呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id: tSimTimerCntlAdapter.cdl 582 2018-12-02 09:20:16Z ertl-hiro $
 */
[singleton, active]
celltype tSimTimerCntlAdapter {
	call	sSimTimerCntl	cSimTimerCntl;
};
