/*
 *		C言語で記述されたアプリケーションから，TECSベースのシリアルイン
 *		タフェースドライバを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id: tSerialAdapter.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */
[singleton, active]
celltype tSerialAdapter {
	call	sSerialPort		cSerialPort[];
};
