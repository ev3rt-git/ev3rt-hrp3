/*
 *		C言語で記述されたアプリケーションから，TECSベースのシステムログ
 *		機能を呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id: tSysLogAdapter.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */
[singleton, active]
celltype tSysLogAdapter {
	call	sSysLog		cSysLog;
};
