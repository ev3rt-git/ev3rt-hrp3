/*
 *		テスト用プラットフォーム（ミューテックス機能の整合性検査付き）
 *		のコンポーネント記述ファイル
 *
 *  $Id: test_pf_bitmutex.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */

/*
 *  テスト用プラットフォームのコンポーネント記述ファイル
 */
import("test_pf.cdl");

/*
 *  ミューテックス機能の整合性検査のセルタイプと組上げ記述
 */
[singleton]
celltype tBitMutex {
	entry	sBuiltInTest	eBuiltInTest;
};

cell tBitMutex BitMutex {					/* テストサービスに接続 */
	eBuiltInTest <= rKernelDomain::TestService.cBuiltInTest;
};
